** Profile: "SCHEMATIC1-yrri"  [ e:\university\electronics 3\lab\6th\sim\gae-schematic1-yrri.sim ] 

** Creating circuit file "gae-schematic1-yrri.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of h:\softwares\orcad\new\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 800ns 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\gae-SCHEMATIC1.net" 


.END
