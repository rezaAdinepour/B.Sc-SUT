** Profile: "SCHEMATIC1-hg"  [ E:\University\Communication Circuits\LAB\5\az5-SCHEMATIC1-hg.sim ] 

** Creating circuit file "az5-SCHEMATIC1-hg.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of h:\softwares\orcad\new\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\az5-SCHEMATIC1.net" 


.END
