** Profile: "SCHEMATIC1-wefe"  [ e:\university\communication circuits\lab\6\az6-schematic1-wefe.sim ] 

** Creating circuit file "az6-schematic1-wefe.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of h:\softwares\orcad\new\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 5��m�s 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\az6-SCHEMATIC1.net" 


.END
