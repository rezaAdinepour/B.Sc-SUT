** Profile: "SCHEMATIC1-Pulse_HW01"  [ E:\UNIVERSITY\ELECTERICAL\Pulse Technique\Dr Ahmadifard\HW\HW01\Simulation\pulse_hw01-SCHEMATIC1-Pulse_HW01.sim ] 

** Creating circuit file "pulse_hw01-SCHEMATIC1-Pulse_HW01.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 20ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pulse_hw01-SCHEMATIC1.net" 


.END
