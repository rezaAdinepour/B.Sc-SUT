** Profile: "SCHEMATIC1-Pulse-HW01"  [ d:\drive e\university\ta\pulse technique\dr ahmadifard\spring 01-02\hws\hw01\simulation\pulse-hw01-schematic1-pulse-hw01.sim ] 

** Creating circuit file "pulse-hw01-schematic1-pulse-hw01.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10us 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pulse-hw01-SCHEMATIC1.net" 


.END
