** Profile: "SCHEMATIC1-Pulse_HW06"  [ E:\UNIVERSITY\ELECTERICAL\PULSE TECHNIQUE\DR AHMADIFARD\SPRING 00-01\HW\HW06\Simulation\8-12\pulse_hw06-SCHEMATIC1-Pulse_HW06.sim ] 

** Creating circuit file "pulse_hw06-SCHEMATIC1-Pulse_HW06.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 200us 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pulse_hw06-SCHEMATIC1.net" 


.END
