** Profile: "SCHEMATIC1-h"  [ E:\UNIVERSITY\Electronics 2\LAB\3rd\currentmirror-SCHEMATIC1-h.sim ] 

** Creating circuit file "currentmirror-SCHEMATIC1-h.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of h:\softwares\orcad\new\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10 10 1gig
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\currentmirror-SCHEMATIC1.net" 


.END
