** Profile: "SCHEMATIC1-Elec1_Lab3"  [ E:\UNIVERSITY\ELECTERICAL\LABS\ELECTRONICS 1\REPORTS\Lab3\Simulation\elec1_lab3-SCHEMATIC1-Elec1_Lab3.sim ] 

** Creating circuit file "elec1_lab3-SCHEMATIC1-Elec1_Lab3.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 3ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\elec1_lab3-SCHEMATIC1.net" 


.END
