** Profile: "SCHEMATIC1-jhu"  [ E:\UNIVERSITY\ELECTRONICS 2\LAB\2ND\SIM\cascodeamp-SCHEMATIC1-jhu.sim ] 

** Creating circuit file "cascodeamp-SCHEMATIC1-jhu.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of h:\softwares\orcad\new\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.4ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\cascodeamp-SCHEMATIC1.net" 


.END
