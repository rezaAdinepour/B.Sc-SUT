** Profile: "SCHEMATIC1-Elec1_Lab8"  [ e:\university\electerical\labs\electronics 1\reports\lab8\simulation\elec1_lab8-schematic1-elec1_lab8.sim ] 

** Creating circuit file "elec1_lab8-schematic1-elec1_lab8.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 5ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\elec1_lab8-SCHEMATIC1.net" 


.END
