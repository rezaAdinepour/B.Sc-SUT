** Profile: "SCHEMATIC1-hj"  [ E:\UNIVERSITY\Electronics 2\LAB\4th\Sim\xff-SCHEMATIC1-hj.sim ] 

** Creating circuit file "xff-SCHEMATIC1-hj.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of h:\softwares\orcad\new\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10 1 100gig
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\xff-SCHEMATIC1.net" 


.END
