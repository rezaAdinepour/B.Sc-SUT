** Profile: "SCHEMATIC1-Elec1_Lab11"  [ E:\UNIVERSITY\ELECTERICAL\LABS\ELECTRONICS 1\Reports\Lab11\Simulation\elec1_lab11-SCHEMATIC1-Elec1_Lab11.sim ] 

** Creating circuit file "elec1_lab11-SCHEMATIC1-Elec1_Lab11.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 1K 1 1000K
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\elec1_lab11-SCHEMATIC1.net" 


.END
