** Profile: "SCHEMATIC1-dfvvs"  [ c:\users\reza\desktop\pspice\project7-SCHEMATIC1-dfvvs.sim ] 

** Creating circuit file "project7-SCHEMATIC1-dfvvs.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 5m 1m 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\project7-SCHEMATIC1.net" 


.END
