** Profile: "SCHEMATIC1-kjk"  [ E:\University\Communication Circuits\LAB\3\az3-SCHEMATIC1-kjk.sim ] 

** Creating circuit file "az3-SCHEMATIC1-kjk.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of h:\softwares\orcad\new\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\az3-SCHEMATIC1.net" 


.END
