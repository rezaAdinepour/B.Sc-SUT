** Profile: "SCHEMATIC1-Elec2_Lab4"  [ e:\university\electerical\labs\electronics 1\reports\lab4\simulation\elec2_lab4-schematic1-elec2_lab4.sim ] 

** Creating circuit file "elec2_lab4-schematic1-elec2_lab4.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 30m 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\elec2_lab4-SCHEMATIC1.net" 


.END
