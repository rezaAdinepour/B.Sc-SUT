** Profile: "SCHEMATIC1-jhgkl;"  [ e:\university\electronics 3\lab\8th\sim\jryk-schematic1-jhgkl;.sim ] 

** Creating circuit file "jryk-schematic1-jhgkl;.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of h:\softwares\orcad\new\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 20s 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\jryk-SCHEMATIC1.net" 


.END
