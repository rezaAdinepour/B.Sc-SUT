** Profile: "SCHEMATIC1-Pulse_HW09"  [ e:\university\electerical\pulse technique\dr ahmadifard\spring 00-01\hw\hw09\simulation\pulse-hw09-schematic1-pulse_hw09.sim ] 

** Creating circuit file "pulse-hw09-schematic1-pulse_hw09.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 40ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pulse-hw09-SCHEMATIC1.net" 


.END
