** Profile: "SCHEMATIC1-Pulse_HW07_Q36"  [ E:\UNIVERSITY\ELECTERICAL\PULSE TECHNIQUE\DR AHMADIFARD\SPRING 00-01\HW\HW07\SIMULATION\Q32\pulse_hw07_q36-SCHEMATIC1-Pulse_HW07_Q36.sim ] 

** Creating circuit file "pulse_hw07_q36-SCHEMATIC1-Pulse_HW07_Q36.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 20ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pulse_hw07_q36-SCHEMATIC1.net" 


.END
