** Profile: "SCHEMATIC1-Elec1_Lab5"  [ E:\UNIVERSITY\ELECTERICAL\LABS\ELECTRONICS 1\REPORTS\LAB5\elec1_lab5-SCHEMATIC1-Elec1_Lab5.sim ] 

** Creating circuit file "elec1_lab5-SCHEMATIC1-Elec1_Lab5.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\elec1_lab5-SCHEMATIC1.net" 


.END
