** Profile: "SCHEMATIC1-Elec1_Lab7"  [ E:\UNIVERSITY\ELECTERICAL\LABS\ELECTRONICS 1\REPORTS\LAB7\SIMULATION\elec1_lab7-SCHEMATIC1-Elec1_Lab7.sim ] 

** Creating circuit file "elec1_lab7-SCHEMATIC1-Elec1_Lab7.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 20ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\elec1_lab7-SCHEMATIC1.net" 


.END
