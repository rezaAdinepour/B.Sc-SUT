** Profile: "SCHEMATIC1-Elec1_Lab2"  [ e:\university\electerical\labs\electronics 1\reports\lab2\simulation\elec1_lab2-schematic1-elec1_lab2.sim ] 

** Creating circuit file "elec1_lab2-schematic1-elec1_lab2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\elec1_lab2-SCHEMATIC1.net" 


.END
