** Profile: "SCHEMATIC1-egrg"  [ E:\UNIVERSITY\Electronics 2\LAB\6th\Sim\gui-SCHEMATIC1-egrg.sim ] 

** Creating circuit file "gui-SCHEMATIC1-egrg.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of h:\softwares\orcad\new\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10 1 100gig
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\gui-SCHEMATIC1.net" 


.END
