** Profile: "SCHEMATIC1-Elec1Lab_Final"  [ E:\UNIVERSITY\ELECTERICAL\LABS\ELECTRONICS 1\Reports\Finall\Simulation\elec1lab_finall-SCHEMATIC1-Elec1Lab_Final.sim ] 

** Creating circuit file "elec1lab_finall-SCHEMATIC1-Elec1Lab_Final.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 1K 1 1000K
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\elec1lab_finall-SCHEMATIC1.net" 


.END
