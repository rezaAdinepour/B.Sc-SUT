** Profile: "SCHEMATIC1-s"  [ e:\university\electronics 3\lab\2nd\sim\diffamp-schematic1-s.sim ] 

** Creating circuit file "diffamp-schematic1-s.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of h:\softwares\orcad\new\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10 10 100gig
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\diffamp-SCHEMATIC1.net" 


.END
