** Profile: "SCHEMATIC1-try1"  [ c:\users\reza\desktop\pspice\project7-schematic1-try1.sim ] 

** Creating circuit file "project7-schematic1-try1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 8m 0 100n 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\project7-SCHEMATIC1.net" 


.END
