** Profile: "SCHEMATIC1-E1_Lab1"  [ e:\university\electerical\labs\electronics 1\reports\lab1\simulation\e1_lab1-schematic1-e1_lab1.sim ] 

** Creating circuit file "e1_lab1-schematic1-e1_lab1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\e1_lab1-SCHEMATIC1.net" 


.END
