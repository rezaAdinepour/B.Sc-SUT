** Profile: "SCHEMATIC1-try2"  [ c:\users\reza\desktop\pspice\project7-SCHEMATIC1-try2.sim ] 

** Creating circuit file "project7-SCHEMATIC1-try2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\project7-SCHEMATIC1.net" 


.END
