** Profile: "SCHEMATIC1-Elec1_Lab6"  [ e:\university\electerical\labs\electronics 1\reports\lab6\simulation\elec1_lab6-schematic1-elec1_lab6.sim ] 

** Creating circuit file "elec1_lab6-schematic1-elec1_lab6.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 20m 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\elec1_lab6-SCHEMATIC1.net" 


.END
