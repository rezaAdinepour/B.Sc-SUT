** Profile: "SCHEMATIC1-vr"  [ e:\university\electronics 3\lab\5th\sim\gwg-schematic1-vr.sim ] 

** Creating circuit file "gwg-schematic1-vr.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of h:\softwares\orcad\new\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 20ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\gwg-SCHEMATIC1.net" 


.END
